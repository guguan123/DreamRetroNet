  D � � � 6Det gick inte att öppna URL %0U i inbyggd webbläsare ;Det gick inte att starta Ovi Webbläsare för webb­program Nej >Inga webb­program är angivna för det här start­programmet COvi Webbläsare hittades inte i din telefon. Ladda ned från Butik? Ja